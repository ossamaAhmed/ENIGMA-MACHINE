library IEEE;
use ieee.std_logic_1164.all;

entity g22_permutation is
port(
	 input_code : in std_logic_vector(4 downto 0);
	 rotor_type : in std_logic_vector(1 downto 0);
	 output_code : out std_logic_vector(4 downto 0);
	 inv_output_code : out std_logic_vector(4 downto 0));
end g22_permutation;

architecture g22_permutation_behavior of g22_permutation is

begin
process (input_code, rotor_type)
begin
   -- Rotor Number One
	if rotor_type = "00" then
			case input_code is
				when "00000" =>
					output_code <=  "00100";
					inv_output_code <=  "10100";
				when "00001" =>
					output_code <=  "01010";
					inv_output_code <=  "10110";
				when  "00010" =>
					output_code <=  "01100";
					inv_output_code <= "11000";
				when  "00011" =>
					output_code <=  "00101";
					inv_output_code <=  "00110";
				when  "00100" =>
					output_code <=  "01011";
					inv_output_code <= "00000";
				when  "00101" =>
					output_code <=  "00110";
					inv_output_code <=  "00011";
				when  "00110" =>
					output_code <=  "00011";
					inv_output_code <=  "00101";
				when  "00111" =>
					output_code <=  "10000";
					inv_output_code <=  "01111";
				when  "01000" =>
					output_code <=  "10101";
					inv_output_code <=  "10101";
				when  "01001" =>
					output_code <= "11001";
					inv_output_code <= "11001";
				when  "01010" =>
					output_code <=  "01101";
					inv_output_code <= "00001";
				when  "01011" =>
					output_code <=  "10011";
					inv_output_code <=  "00100";
				when  "01100" =>
					output_code <=  "01110";
					inv_output_code <=  "00010";
				when  "01101" =>
					output_code <=  "10110";
					inv_output_code <=  "01010";
				when  "01110" =>
					output_code <= "11000";
					inv_output_code <=  "01100";
				when  "01111" =>
					output_code <=  "00111";
					inv_output_code <=  "10011";
				when  "10000" =>
					output_code <= "10111";
					inv_output_code <=  "00111";
				when  "10001" =>
					output_code <=  "10100";
					inv_output_code <= "10111";
				when  "10010" =>
					output_code <=  "10010";
					inv_output_code <=  "10010";
				when  "10011" =>
					output_code <=  "01111";
					inv_output_code <=  "01011";
				when  "10100" =>
					output_code <= "00000";
					inv_output_code <=  "10001";
				when  "10101" =>
					output_code <=  "01000";
					inv_output_code <=  "01000";
				when  "10110" =>
					output_code <= "00001";
					inv_output_code <=  "01101";
				when "10111" =>
					output_code <=  "10001";
					inv_output_code <=  "10000";
				when "11000" =>
					output_code <=  "00010";
					inv_output_code <=  "01110";
				when "11001" =>
					output_code <=  "01001";
					inv_output_code <=  "01001";
				when others =>
					output_code <= "11111";
					inv_output_code <= "11111";
			end case;
			-- Rotor Number two
		elsif rotor_type = "01" then
			case input_code is
				when "00000" =>
					output_code <= "00000";
					inv_output_code <= "00000";
				when "00001" =>
					output_code <=  "01001";
					inv_output_code <=  "01001";
				when  "00010" =>
					output_code <=  "00011";
					inv_output_code <=  "01111";
				when  "00011" =>
					output_code <=  "01010";
					inv_output_code <=  "00010";
				when  "00100" =>
					output_code <=  "10010";
					inv_output_code <= "11001";
				when  "00101" =>
					output_code <=  "01000";
					inv_output_code <=  "10110";
				when  "00110" =>
					output_code <=  "10001";
					inv_output_code <=  "10001";
				when  "00111" =>
					output_code <=  "10100";
					inv_output_code <=  "01011";
				when  "01000" =>
					output_code <= "10111";
					inv_output_code <=  "00101";
				when  "01001" =>
					output_code <= "00001";
					inv_output_code <= "00001";
				when  "01010" =>
					output_code <=  "01011";
					inv_output_code <=  "00011";
				when  "01011" =>
					output_code <=  "00111";
					inv_output_code <=  "01010";
				when  "01100" =>
					output_code <=  "10110";
					inv_output_code <=  "01110";
				when  "01101" =>
					output_code <=  "10011";
					inv_output_code <=  "10011";
				when  "01110" =>
					output_code <=  "01100";
					inv_output_code <= "11000";
				when  "01111" =>
					output_code <=  "00010";
					inv_output_code <=  "10100";
				when  "10000" =>
					output_code <=  "10000";
					inv_output_code <=  "10000";
				when  "10001" =>
					output_code <=  "00110";
					inv_output_code <=  "00110";
				when  "10010" =>
					output_code <= "11001";
					inv_output_code <=  "00100";
				when  "10011" =>
					output_code <=  "01101";
					inv_output_code <=  "01101";
				when  "10100" =>
					output_code <=  "01111";
					inv_output_code <=  "00111";
				when  "10101" =>
					output_code <= "11000";
					inv_output_code <= "10111";
				when  "10110" =>
					output_code <=  "00101";
					inv_output_code <=  "01100";
				when "10111" =>
					output_code <=  "10101";
					inv_output_code <=  "01000";
				when "11000" =>
					output_code <=  "01110";
					inv_output_code <=  "10101";
				when "11001" =>
					output_code <=  "00100";
					inv_output_code <=  "10010";
				when others =>
					output_code <= "11111";
					inv_output_code <= "11111";
			end case;
			-- Rotor Number Three
		elsif rotor_type = "10" then
			case input_code is
				when "00000" =>
					output_code <= "00001";
					inv_output_code <=  "10011";
				when "00001" =>
					output_code <=  "00011";
					inv_output_code <= "00000";
				when  "00010" =>
					output_code <=  "00101";
					inv_output_code <=  "00110";
				when  "00011" =>
					output_code <=  "00111";
					inv_output_code <=  "00011";
				when  "00100" =>
					output_code <=  "01001";
					inv_output_code <=  "01111";
				when  "00101" =>
					output_code <=  "01011";
					inv_output_code <=  "00010";
				when  "00110" =>
					output_code <=  "00010";
					inv_output_code <=  "10010";
				when  "00111" =>
					output_code <=  "01111";
					inv_output_code <=  "00011";
				when  "01000" =>
					output_code <=  "10001";
					inv_output_code <=  "10000";
				when  "01001" =>
					output_code <=  "10011";
					inv_output_code <=  "00100";
				when  "01010" =>
					output_code <= "10111";
					inv_output_code <=  "10100";
				when  "01011" =>
					output_code <=  "10101";
					inv_output_code <=  "00101";
				when  "01100" =>
					output_code <= "11001";
					inv_output_code <=  "10101";
				when  "01101" =>
					output_code <=  "01101";
					inv_output_code <=  "01101";
				when  "01110" =>
					output_code <= "11000";
					inv_output_code <= "11001";
				when  "01111" =>
					output_code <=  "00100";
					inv_output_code <=  "00111";
				when  "10000" =>
					output_code <=  "01000";
					inv_output_code <= "11000";
				when  "10001" =>
					output_code <=  "10110";
					inv_output_code <=  "01000";
				when  "10010" =>
					output_code <=  "00110";
					inv_output_code <= "10111";
				when  "10011" =>
					output_code <= "00000";
					inv_output_code <=  "01001";
				when  "10100" =>
					output_code <=  "01010";
					inv_output_code <=  "10110";
				when  "10101" =>
					output_code <=  "01100";
					inv_output_code <=  "01011";
				when  "10110" =>
					output_code <=  "10100";
					inv_output_code <=  "10001";
				when "10111" =>
					output_code <=  "10010";
					inv_output_code <=  "01010";
				when "11000" =>
					output_code <=  "10000";
					inv_output_code <=  "01110";
				when "11001" =>
					output_code <=  "01110";
					inv_output_code <=  "01100";
				when others =>
					output_code <= "11111";
					inv_output_code <= "11111";
				end case;			
		-- Rotor Number Four  
		elsif rotor_type = "11" then
			case input_code is
				when "00000" =>
					output_code <=  "00100";
					inv_output_code <=  "00111";
				when "00001" =>
					output_code <=  "10010";
					inv_output_code <= "11001";
				when  "00010" =>
					output_code <=  "01110";
					inv_output_code <=  "10110";
				when  "00011" =>
					output_code <=  "10101";
					inv_output_code <=  "10101";
				when  "00100" =>
					output_code <=  "01111";
					inv_output_code <= "00000";
				when  "00101" =>
					output_code <= "11001";
					inv_output_code <=  "10001";
				when  "00110" =>
					output_code <=  "01001";
					inv_output_code <=  "10011";
				when  "00111" =>
					output_code <= "00000";
					inv_output_code <=  "01101";
				when  "01000" =>
					output_code <= "11000";
					inv_output_code <=  "01011";
				when  "01001" =>
					output_code <=  "10000";
					inv_output_code <=  "00110";
				when  "01010" =>
					output_code <=  "10100";
					inv_output_code <=  "10100";
				when  "01011" =>
					output_code <=  "01000";
					inv_output_code <=  "01111";
				when  "01100" =>
					output_code <=  "10001";
					inv_output_code <= "10111";
				when  "01101" =>
					output_code <=  "00111";
					inv_output_code <=  "10000";
				when  "01110" =>
					output_code <= "10111";
					inv_output_code <=  "00010";
				when  "01111" =>
					output_code <=  "01011";
					inv_output_code <=  "00100";
				when  "10000" =>
					output_code <=  "01101";
					inv_output_code <=  "01001";
				when  "10001" =>
					output_code <=  "00101";
					inv_output_code <=  "01100";
				when  "10010" =>
					output_code <=  "10011";
					inv_output_code <= "00001";
				when  "10011" =>
					output_code <=  "00110";
					inv_output_code <=  "10010";
				when  "10100" =>
					output_code <=  "01010";
					inv_output_code <=  "01010";
				when  "10101" =>
					output_code <=  "00011";
					inv_output_code <=  "00011";
				when  "10110" =>
					output_code <=  "00010";
					inv_output_code <= "11000";
				when "10111" =>
					output_code <=  "01100";
					inv_output_code <=  "01110";
				when "11000" =>
					output_code <=  "10110";
					inv_output_code <=  "01000";
				when "11001" =>
					output_code <= "00001";
					inv_output_code <=  "00101";
				when others =>
					output_code <= "11111";
					inv_output_code <= "11111";
			end case;
		end if;
end process;

end g22_permutation_behavior;